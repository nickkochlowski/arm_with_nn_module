package fsm_pkg_1;

	typedef enum logic [2:0] {s0 = 3'b000, 
				s1 = 3'b001, 
				s2 = 3'b010,
				s3 = 3'b011,
				s4 = 3'b100, 
				  XX = 3'bxxx} state_1;
endpackage
