package fsm_pkg_2;

	typedef enum logic [4:0] {s0 = 5'b00000,
				s1 = 5'b00001, 
				s2 = 5'b00010,
				s3 = 5'b00011,
				s4 = 5'b00100, 
				s5 = 5'b00101, 
				s6 = 5'b00110, 
				s7 = 5'b00111, 
				s8 = 5'b01000, 
				s9 = 5'b01001, 
				s10 = 5'b01010, 
				s11 = 5'b01011, 
				s12 = 5'b01100, 
				s13 = 5'b01101, 
				s14 = 5'b01110,
				s15 = 5'b01111,
				s16 = 5'b10000,
				XX = 5'bxxxxx} state_2;
endpackage
